module Not (input a, output res);
    C1 C (1'b1, 1'b0, a, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, res);
endmodule