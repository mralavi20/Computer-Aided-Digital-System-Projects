module Adder (input [7:0] data_in1, data_in2, output [7:0] data_out);
    assign data_out = data_in1 + data_in2;
endmodule