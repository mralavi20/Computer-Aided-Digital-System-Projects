module And (input a, b, output res);
    C1 C (1'b0, b, a, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, res);
endmodule