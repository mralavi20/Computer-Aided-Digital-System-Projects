module Nand (input a, b, output res);
    C1 C (1'b1, 1'b1, 1'b1, 1'b1, 1'b0, b, a, 1'b0, res);
endmodule
