module Or (input a, b, output res);
    C1 C (b, 1'b1, a, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, res);
endmodule